/*

Copyright (c) 2017 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * FPGA top-level module
 */
module fpga (
    /*
     * Clock: 125MHz LVDS
     * Reset: Push button, active low
     */
    input  wire       clk_125mhz_p,
    input  wire       clk_125mhz_n,
    input  wire       reset,

    /*
     * GPIO
     */
    input  wire       btnu,
    input  wire       btnl,
    input  wire       btnd,
    input  wire       btnr,
    input  wire       btnc,
    input  wire [3:0] sw,
    output wire [7:0] led,

    /*
     * I2C for board management
     */
    inout  wire       i2c_scl,
    inout  wire       i2c_sda,

    /*
     * Ethernet: QSFP28
     */
    output wire       qsfp1_tx1_p,
    output wire       qsfp1_tx1_n,
    input  wire       qsfp1_rx1_p,
    input  wire       qsfp1_rx1_n,
    output wire       qsfp1_tx2_p,
    output wire       qsfp1_tx2_n,
    input  wire       qsfp1_rx2_p,
    input  wire       qsfp1_rx2_n,
    output wire       qsfp1_tx3_p,
    output wire       qsfp1_tx3_n,
    input  wire       qsfp1_rx3_p,
    input  wire       qsfp1_rx3_n,
    output wire       qsfp1_tx4_p,
    output wire       qsfp1_tx4_n,
    input  wire       qsfp1_rx4_p,
    input  wire       qsfp1_rx4_n,
    input  wire       qsfp1_mgt_refclk_0_p,
    input  wire       qsfp1_mgt_refclk_0_n,
    // input  wire       qsfp1_mgt_refclk_1_p,
    // input  wire       qsfp1_mgt_refclk_1_n,
    // output wire       qsfp1_recclk_p,
    // output wire       qsfp1_recclk_n,
    output wire       qsfp1_modsell,
    output wire       qsfp1_resetl,
    input  wire       qsfp1_modprsl,
    input  wire       qsfp1_intl,
    output wire       qsfp1_lpmode,

    output wire       qsfp2_tx1_p,
    output wire       qsfp2_tx1_n,
    input  wire       qsfp2_rx1_p,
    input  wire       qsfp2_rx1_n,
    output wire       qsfp2_tx2_p,
    output wire       qsfp2_tx2_n,
    input  wire       qsfp2_rx2_p,
    input  wire       qsfp2_rx2_n,
    output wire       qsfp2_tx3_p,
    output wire       qsfp2_tx3_n,
    input  wire       qsfp2_rx3_p,
    input  wire       qsfp2_rx3_n,
    output wire       qsfp2_tx4_p,
    output wire       qsfp2_tx4_n,
    input  wire       qsfp2_rx4_p,
    input  wire       qsfp2_rx4_n,
    // input  wire       qsfp2_mgt_refclk_0_p,
    // input  wire       qsfp2_mgt_refclk_0_n,
    // input  wire       qsfp2_mgt_refclk_1_p,
    // input  wire       qsfp2_mgt_refclk_1_n,
    // output wire       qsfp2_recclk_p,
    // output wire       qsfp2_recclk_n,
    output wire       qsfp2_modsell,
    output wire       qsfp2_resetl,
    input  wire       qsfp2_modprsl,
    input  wire       qsfp2_intl,
    output wire       qsfp2_lpmode,

    /*
     * Ethernet: 1000BASE-T SGMII
     */
    input  wire       phy_sgmii_rx_p,
    input  wire       phy_sgmii_rx_n,
    output wire       phy_sgmii_tx_p,
    output wire       phy_sgmii_tx_n,
    input  wire       phy_sgmii_clk_p,
    input  wire       phy_sgmii_clk_n,
    output wire       phy_reset_n,
    input  wire       phy_int_n,
    inout  wire       phy_mdio,
    output wire       phy_mdc,

    /*
     * UART: 115200 bps, 8N1
     */
    input  wire       uart_rxd,
    output wire       uart_txd,
    output wire       uart_rts,
    input  wire       uart_cts
);

// Clock and reset

wire clk_125mhz_ibufg;
wire clk_125mhz_mmcm_out;
wire clk_62mhz_mmcm_out;

// Internal 125 MHz clock
wire clk_125mhz_int;
wire rst_125mhz_int;

// Internal 62.5 MHz clock
wire clk_62mhz_int;
wire rst_62mhz_int;

wire mmcm_rst = reset;
wire mmcm_locked;
wire mmcm_clkfb;

IBUFGDS #(
   .DIFF_TERM("FALSE"),
   .IBUF_LOW_PWR("FALSE")   
)
clk_125mhz_ibufg_inst (
   .O   (clk_125mhz_ibufg),
   .I   (clk_125mhz_p),
   .IB  (clk_125mhz_n) 
);

// MMCM instance
// 125 MHz in, 125 MHz out
// PFD range: 10 MHz to 500 MHz
// VCO range: 800 MHz to 1600 MHz
// M = 8, D = 1 sets Fvco = 1000 MHz (in range)
// Divide by 8 to get output frequency of 125 MHz
// Divide by 16 to get output frequency of 62.5 MHz
MMCME4_BASE #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKOUT0_DIVIDE_F(8),
    .CLKOUT0_DUTY_CYCLE(0.5),
    .CLKOUT0_PHASE(0),
    .CLKOUT1_DIVIDE(16),
    .CLKOUT1_DUTY_CYCLE(0.5),
    .CLKOUT1_PHASE(0),
    .CLKOUT2_DIVIDE(1),
    .CLKOUT2_DUTY_CYCLE(0.5),
    .CLKOUT2_PHASE(0),
    .CLKOUT3_DIVIDE(1),
    .CLKOUT3_DUTY_CYCLE(0.5),
    .CLKOUT3_PHASE(0),
    .CLKOUT4_DIVIDE(1),
    .CLKOUT4_DUTY_CYCLE(0.5),
    .CLKOUT4_PHASE(0),
    .CLKOUT5_DIVIDE(1),
    .CLKOUT5_DUTY_CYCLE(0.5),
    .CLKOUT5_PHASE(0),
    .CLKOUT6_DIVIDE(1),
    .CLKOUT6_DUTY_CYCLE(0.5),
    .CLKOUT6_PHASE(0),
    .CLKFBOUT_MULT_F(8),
    .CLKFBOUT_PHASE(0),
    .DIVCLK_DIVIDE(1),
    .REF_JITTER1(0.010),
    .CLKIN1_PERIOD(8.0),
    .STARTUP_WAIT("FALSE"),
    .CLKOUT4_CASCADE("FALSE")
)
clk_mmcm_inst (
    .CLKIN1(clk_125mhz_ibufg),
    .CLKFBIN(mmcm_clkfb),
    .RST(mmcm_rst),
    .PWRDWN(1'b0),
    .CLKOUT0(clk_125mhz_mmcm_out),
    .CLKOUT0B(),
    .CLKOUT1(clk_62mhz_mmcm_out),
    .CLKOUT1B(),
    .CLKOUT2(),
    .CLKOUT2B(),
    .CLKOUT3(),
    .CLKOUT3B(),
    .CLKOUT4(),
    .CLKOUT5(),
    .CLKOUT6(),
    .CLKFBOUT(mmcm_clkfb),
    .CLKFBOUTB(),
    .LOCKED(mmcm_locked)
);

BUFG
clk_125mhz_bufg_inst (
    .I(clk_125mhz_mmcm_out),
    .O(clk_125mhz_int)
);

BUFG
clk_62mhz_bufg_inst (
    .I(clk_62mhz_mmcm_out),
    .O(clk_62mhz_int)
);

sync_reset #(
    .N(4)
)
sync_reset_125mhz_inst (
    .clk(clk_125mhz_int),
    .rst(~mmcm_locked),
    .out(rst_125mhz_int)
);

sync_reset #(
    .N(4)
)
sync_reset_62mhz_inst (
    .clk(clk_62mhz_int),
    .rst(~mmcm_locked),
    .out(rst_62mhz_int)
);

// GPIO
wire btnu_int;
wire btnl_int;
wire btnd_int;
wire btnr_int;
wire btnc_int;
wire [3:0] sw_int;

debounce_switch #(
    .WIDTH(9),
    .N(4),
    .RATE(125000)
)
debounce_switch_inst (
    .clk(clk_125mhz_int),
    .rst(rst_125mhz_int),
    .in({btnu,
        btnl,
        btnd,
        btnr,
        btnc,
        sw}),
    .out({btnu_int,
        btnl_int,
        btnd_int,
        btnr_int,
        btnc_int,
        sw_int})
);

wire uart_rxd_int;
wire uart_cts_int;

sync_signal #(
    .WIDTH(2),
    .N(2)
)
sync_signal_inst (
    .clk(clk_125mhz_int),
    .in({uart_rxd, uart_cts}),
    .out({uart_rxd_int, uart_cts_int})
);

wire i2c_scl_i;
wire i2c_scl_o;
wire i2c_scl_t;
wire i2c_sda_i;
wire i2c_sda_o;
wire i2c_sda_t;

assign i2c_scl_i = i2c_scl;
assign i2c_scl = i2c_scl_t ? 1'bz : i2c_scl_o;
assign i2c_sda_i = i2c_sda;
assign i2c_sda = i2c_sda_t ? 1'bz : i2c_sda_o;

// GTY instances
assign qsfp1_modsell = 1'b0;
assign qsfp1_resetl = 1'b1;
assign qsfp1_lpmode = 1'b0;

assign qsfp2_modsell = 1'b0;
assign qsfp2_resetl = 1'b1;
assign qsfp2_lpmode = 1'b0;

wire gty_drp_clk = clk_62mhz_int;
wire gty_drp_rst = rst_62mhz_int;

wire [7:0] xfcp_mgt_up_tdata;
wire xfcp_mgt_up_tvalid;
wire xfcp_mgt_up_tready;
wire xfcp_mgt_up_tlast;
wire xfcp_mgt_up_tuser;
wire [7:0] xfcp_mgt_down_tdata;
wire xfcp_mgt_down_tvalid;
wire xfcp_mgt_down_tready;
wire xfcp_mgt_down_tlast;
wire xfcp_mgt_down_tuser;

wire [7:0] xfcp_mgt_fifo_up_tdata;
wire xfcp_mgt_fifo_up_tvalid;
wire xfcp_mgt_fifo_up_tready;
wire xfcp_mgt_fifo_up_tlast;
wire xfcp_mgt_fifo_up_tuser;
wire [7:0] xfcp_mgt_fifo_down_tdata;
wire xfcp_mgt_fifo_down_tvalid;
wire xfcp_mgt_fifo_down_tready;
wire xfcp_mgt_fifo_down_tlast;
wire xfcp_mgt_fifo_down_tuser;

wire [7:0] xfcp_qsfp1_gty_up_tdata;
wire xfcp_qsfp1_gty_up_tvalid;
wire xfcp_qsfp1_gty_up_tready;
wire xfcp_qsfp1_gty_up_tlast;
wire xfcp_qsfp1_gty_up_tuser;
wire [7:0] xfcp_qsfp1_gty_down_tdata;
wire xfcp_qsfp1_gty_down_tvalid;
wire xfcp_qsfp1_gty_down_tready;
wire xfcp_qsfp1_gty_down_tlast;
wire xfcp_qsfp1_gty_down_tuser;

wire [7:0] xfcp_qsfp2_gty_up_tdata;
wire xfcp_qsfp2_gty_up_tvalid;
wire xfcp_qsfp2_gty_up_tready;
wire xfcp_qsfp2_gty_up_tlast;
wire xfcp_qsfp2_gty_up_tuser;
wire [7:0] xfcp_qsfp2_gty_down_tdata;
wire xfcp_qsfp2_gty_down_tvalid;
wire xfcp_qsfp2_gty_down_tready;
wire xfcp_qsfp2_gty_down_tlast;
wire xfcp_qsfp2_gty_down_tuser;

axis_async_fifo #(
    .DEPTH(32),
    .DATA_WIDTH(8)
)
xfcp_mgt_fifo_down (
    // Common reset
    .async_rst(rst_125mhz_int | gty_drp_rst),
    // AXI input
    .s_clk(clk_125mhz_int),
    .s_axis_tdata(xfcp_mgt_down_tdata),
    .s_axis_tvalid(xfcp_mgt_down_tvalid),
    .s_axis_tready(xfcp_mgt_down_tready),
    .s_axis_tlast(xfcp_mgt_down_tlast),
    .s_axis_tuser(xfcp_mgt_down_tuser),
    // AXI output
    .m_clk(gty_drp_clk),
    .m_axis_tdata(xfcp_mgt_fifo_down_tdata),
    .m_axis_tvalid(xfcp_mgt_fifo_down_tvalid),
    .m_axis_tready(xfcp_mgt_fifo_down_tready),
    .m_axis_tlast(xfcp_mgt_fifo_down_tlast),
    .m_axis_tuser(xfcp_mgt_fifo_down_tuser)
);

axis_async_fifo #(
    .DEPTH(32),
    .DATA_WIDTH(8)
)
xfcp_mgt_fifo_up (
    // Common reset
    .async_rst(rst_125mhz_int | gty_drp_rst),
    // AXI input
    .s_clk(gty_drp_clk),
    .s_axis_tdata(xfcp_mgt_fifo_up_tdata),
    .s_axis_tvalid(xfcp_mgt_fifo_up_tvalid),
    .s_axis_tready(xfcp_mgt_fifo_up_tready),
    .s_axis_tlast(xfcp_mgt_fifo_up_tlast),
    .s_axis_tuser(xfcp_mgt_fifo_up_tuser),
    // AXI output
    .m_clk(clk_125mhz_int),
    .m_axis_tdata(xfcp_mgt_up_tdata),
    .m_axis_tvalid(xfcp_mgt_up_tvalid),
    .m_axis_tready(xfcp_mgt_up_tready),
    .m_axis_tlast(xfcp_mgt_up_tlast),
    .m_axis_tuser(xfcp_mgt_up_tuser)
);

xfcp_switch #(
    .PORTS(2),
    .XFCP_ID_TYPE(16'h0100),
    .XFCP_ID_STR("XFCP switch"),
    .XFCP_EXT_ID(0),
    .XFCP_EXT_ID_STR("GTY QUADs")
)
xfcp_switch_inst (
    .clk(gty_drp_clk),
    .rst(gty_drp_rst),
    .up_xfcp_in_tdata(xfcp_mgt_fifo_down_tdata),
    .up_xfcp_in_tvalid(xfcp_mgt_fifo_down_tvalid),
    .up_xfcp_in_tready(xfcp_mgt_fifo_down_tready),
    .up_xfcp_in_tlast(xfcp_mgt_fifo_down_tlast),
    .up_xfcp_in_tuser(xfcp_mgt_fifo_down_tuser),
    .up_xfcp_out_tdata(xfcp_mgt_fifo_up_tdata),
    .up_xfcp_out_tvalid(xfcp_mgt_fifo_up_tvalid),
    .up_xfcp_out_tready(xfcp_mgt_fifo_up_tready),
    .up_xfcp_out_tlast(xfcp_mgt_fifo_up_tlast),
    .up_xfcp_out_tuser(xfcp_mgt_fifo_up_tuser),
    .down_xfcp_in_tdata(  {xfcp_qsfp2_gty_up_tdata,    xfcp_qsfp1_gty_up_tdata   }),
    .down_xfcp_in_tvalid( {xfcp_qsfp2_gty_up_tvalid,   xfcp_qsfp1_gty_up_tvalid  }),
    .down_xfcp_in_tready( {xfcp_qsfp2_gty_up_tready,   xfcp_qsfp1_gty_up_tready  }),
    .down_xfcp_in_tlast(  {xfcp_qsfp2_gty_up_tlast,    xfcp_qsfp1_gty_up_tlast   }),
    .down_xfcp_in_tuser(  {xfcp_qsfp2_gty_up_tuser,    xfcp_qsfp1_gty_up_tuser   }),
    .down_xfcp_out_tdata( {xfcp_qsfp2_gty_down_tdata,  xfcp_qsfp1_gty_down_tdata }),
    .down_xfcp_out_tvalid({xfcp_qsfp2_gty_down_tvalid, xfcp_qsfp1_gty_down_tvalid}),
    .down_xfcp_out_tready({xfcp_qsfp2_gty_down_tready, xfcp_qsfp1_gty_down_tready}),
    .down_xfcp_out_tlast( {xfcp_qsfp2_gty_down_tlast,  xfcp_qsfp1_gty_down_tlast }),
    .down_xfcp_out_tuser( {xfcp_qsfp2_gty_down_tuser,  xfcp_qsfp1_gty_down_tuser })
);

// QSFP GTY
assign qsfp1_modsell = 1'b0;
assign qsfp1_resetl = 1'b1;
assign qsfp1_lpmode = 1'b0;

assign qsfp2_modsell = 1'b0;
assign qsfp2_resetl = 1'b1;
assign qsfp2_lpmode = 1'b0;

wire [2*10-1:0] qsfp_gty_com_drp_addr;
wire [2*16-1:0] qsfp_gty_com_drp_do;
wire [2*16-1:0] qsfp_gty_com_drp_di;
wire [2-1:0] qsfp_gty_com_drp_en;
wire [2-1:0] qsfp_gty_com_drp_we;
wire [2-1:0] qsfp_gty_com_drp_rdy;

wire [8*10-1:0] qsfp_gty_drp_addr;
wire [8*16-1:0] qsfp_gty_drp_do;
wire [8*16-1:0] qsfp_gty_drp_di;
wire [8-1:0] qsfp_gty_drp_en;
wire [8-1:0] qsfp_gty_drp_we;
wire [8-1:0] qsfp_gty_drp_rdy;

wire [8-1:0] qsfp_gty_reset;
wire [8-1:0] qsfp_gty_tx_reset;
wire [8-1:0] qsfp_gty_rx_reset;

wire qsfp_gty_txusrclk2;
wire [8*4-1:0] qsfp_gty_txprbssel;
wire [8-1:0] qsfp_gty_txprbsforceerr;
wire [8-1:0] qsfp_gty_txpolarity;
wire [8-1:0] qsfp_gty_txelecidle;
wire [8-1:0] qsfp_gty_txinhibit;
wire [8*5-1:0] qsfp_gty_txdiffctrl;
wire [8*7-1:0] qsfp_gty_txmaincursor;
wire [8*5-1:0] qsfp_gty_txpostcursor;
wire [8*5-1:0] qsfp_gty_txprecursor;

wire qsfp_gty_rxusrclk2;
wire [8-1:0] qsfp_gty_rxpolarity;
wire [8-1:0] qsfp_gty_rxprbscntreset;
wire [8*4-1:0] qsfp_gty_rxprbssel;
wire [8-1:0] qsfp_gty_rxprbserr;
wire [8-1:0] qsfp_gty_rxprbslocked;

xfcp_gty_quad #(
    .CH(4),
    .SW_XFCP_ID_TYPE(16'h0100),
    .SW_XFCP_ID_STR("GTY QUAD 231"),
    .SW_XFCP_EXT_ID(0),
    .SW_XFCP_EXT_ID_STR("QSFP1 GTY QUAD"),
    .COM_XFCP_ID_TYPE(16'h8A92),
    .COM_XFCP_ID_STR("GTY COM X1Y12"),
    .COM_XFCP_EXT_ID(0),
    .COM_XFCP_EXT_ID_STR("QSFP1 GTY COM"),
    .CH_0_XFCP_ID_TYPE(16'h8A93),
    .CH_0_XFCP_ID_STR("GTY CH0 X1Y48"),
    .CH_0_XFCP_EXT_ID(0),
    .CH_0_XFCP_EXT_ID_STR("QSFP1 CH1"),
    .CH_1_XFCP_ID_TYPE(16'h8A93),
    .CH_1_XFCP_ID_STR("GTY CH1 X1Y49"),
    .CH_1_XFCP_EXT_ID(0),
    .CH_1_XFCP_EXT_ID_STR("QSFP1 CH2"),
    .CH_2_XFCP_ID_TYPE(16'h8A93),
    .CH_2_XFCP_ID_STR("GTY CH2 X1Y50"),
    .CH_2_XFCP_EXT_ID(0),
    .CH_2_XFCP_EXT_ID_STR("QSFP1 CH3"),
    .CH_3_XFCP_ID_TYPE(16'h8A93),
    .CH_3_XFCP_ID_STR("GTY CH3 X1Y51"),
    .CH_3_XFCP_EXT_ID(0),
    .CH_3_XFCP_EXT_ID_STR("QSFP1 CH4"),
    .COM_ADDR_WIDTH(10),
    .CH_ADDR_WIDTH(10)
)
xfcp_qsfp1_gty_quad_inst (
    .clk(gty_drp_clk),
    .rst(gty_drp_rst),

    .up_xfcp_in_tdata(xfcp_qsfp1_gty_down_tdata),
    .up_xfcp_in_tvalid(xfcp_qsfp1_gty_down_tvalid),
    .up_xfcp_in_tready(xfcp_qsfp1_gty_down_tready),
    .up_xfcp_in_tlast(xfcp_qsfp1_gty_down_tlast),
    .up_xfcp_in_tuser(xfcp_qsfp1_gty_down_tuser),
    .up_xfcp_out_tdata(xfcp_qsfp1_gty_up_tdata),
    .up_xfcp_out_tvalid(xfcp_qsfp1_gty_up_tvalid),
    .up_xfcp_out_tready(xfcp_qsfp1_gty_up_tready),
    .up_xfcp_out_tlast(xfcp_qsfp1_gty_up_tlast),
    .up_xfcp_out_tuser(xfcp_qsfp1_gty_up_tuser),

    .gty_com_drp_addr(qsfp_gty_com_drp_addr[0*10 +: 10]),
    .gty_com_drp_do(qsfp_gty_com_drp_do[0*16 +: 16]),
    .gty_com_drp_di(qsfp_gty_com_drp_di[0*16 +: 16]),
    .gty_com_drp_en(qsfp_gty_com_drp_en[0*1 +: 1]),
    .gty_com_drp_we(qsfp_gty_com_drp_we[0*1 +: 1]),
    .gty_com_drp_rdy(qsfp_gty_com_drp_rdy[0*1 +: 1]),

    .gty_drp_addr(qsfp_gty_drp_addr[0*4*10 +: 4*10]),
    .gty_drp_do(qsfp_gty_drp_do[0*4*16 +: 4*16]),
    .gty_drp_di(qsfp_gty_drp_di[0*4*16 +: 4*16]),
    .gty_drp_en(qsfp_gty_drp_en[0*4*1 +: 4*1]),
    .gty_drp_we(qsfp_gty_drp_we[0*4*1 +: 4*1]),
    .gty_drp_rdy(qsfp_gty_drp_rdy[0*4*1 +: 4*1]),

    .gty_reset(qsfp_gty_reset[0*4*1 +: 4*1]),
    .gty_tx_reset(qsfp_gty_tx_reset[0*4*1 +: 4*1]),
    .gty_rx_reset(qsfp_gty_rx_reset[0*4*1 +: 4*1]),

    .gty_txusrclk2({4{qsfp_gty_txusrclk2}}),
    .gty_txprbssel(qsfp_gty_txprbssel[0*4*4 +: 4*4]),
    .gty_txprbsforceerr(qsfp_gty_txprbsforceerr[0*4*1 +: 4*1]),
    .gty_txpolarity(qsfp_gty_txpolarity[0*4*1 +: 4*1]),
    .gty_txelecidle(qsfp_gty_txelecidle[0*4*1 +: 4*1]),
    .gty_txinhibit(qsfp_gty_txinhibit[0*4*1 +: 4*1]),
    .gty_txdiffctrl(qsfp_gty_txdiffctrl[0*4*5 +: 4*5]),
    .gty_txmaincursor(qsfp_gty_txmaincursor[0*4*7 +: 4*7]),
    .gty_txpostcursor(qsfp_gty_txpostcursor[0*4*5 +: 4*5]),
    .gty_txprecursor(qsfp_gty_txprecursor[0*4*5 +: 4*5]),

    .gty_rxusrclk2({4{qsfp_gty_rxusrclk2}}),
    .gty_rxpolarity(qsfp_gty_rxpolarity[0*4*1 +: 4*1]),
    .gty_rxprbscntreset(qsfp_gty_rxprbscntreset[0*4*1 +: 4*1]),
    .gty_rxprbssel(qsfp_gty_rxprbssel[0*4*4 +: 4*4]),
    .gty_rxprbserr(qsfp_gty_rxprbserr[0*4*1 +: 4*1]),
    .gty_rxprbslocked(qsfp_gty_rxprbslocked[0*4*1 +: 4*1])
);

xfcp_gty_quad #(
    .CH(4),
    .SW_XFCP_ID_TYPE(16'h0100),
    .SW_XFCP_ID_STR("GTY QUAD 232"),
    .SW_XFCP_EXT_ID(0),
    .SW_XFCP_EXT_ID_STR("QSFP2 GTY QUAD"),
    .COM_XFCP_ID_TYPE(16'h8A92),
    .COM_XFCP_ID_STR("GTY COM X1Y13"),
    .COM_XFCP_EXT_ID(0),
    .COM_XFCP_EXT_ID_STR("QSFP2 GTY COM"),
    .CH_0_XFCP_ID_TYPE(16'h8A93),
    .CH_0_XFCP_ID_STR("GTY CH0 X1Y52"),
    .CH_0_XFCP_EXT_ID(0),
    .CH_0_XFCP_EXT_ID_STR("QSFP2 CH1"),
    .CH_1_XFCP_ID_TYPE(16'h8A93),
    .CH_1_XFCP_ID_STR("GTY CH1 X1Y53"),
    .CH_1_XFCP_EXT_ID(0),
    .CH_1_XFCP_EXT_ID_STR("QSFP2 CH2"),
    .CH_2_XFCP_ID_TYPE(16'h8A93),
    .CH_2_XFCP_ID_STR("GTY CH2 X1Y54"),
    .CH_2_XFCP_EXT_ID(0),
    .CH_2_XFCP_EXT_ID_STR("QSFP2 CH3"),
    .CH_3_XFCP_ID_TYPE(16'h8A93),
    .CH_3_XFCP_ID_STR("GTY CH3 X1Y55"),
    .CH_3_XFCP_EXT_ID(0),
    .CH_3_XFCP_EXT_ID_STR("QSFP2 CH4"),
    .COM_ADDR_WIDTH(10),
    .CH_ADDR_WIDTH(10)
)
xfcp_qsfp2_gty_quad_inst (
    .clk(gty_drp_clk),
    .rst(gty_drp_rst),

    .up_xfcp_in_tdata(xfcp_qsfp2_gty_down_tdata),
    .up_xfcp_in_tvalid(xfcp_qsfp2_gty_down_tvalid),
    .up_xfcp_in_tready(xfcp_qsfp2_gty_down_tready),
    .up_xfcp_in_tlast(xfcp_qsfp2_gty_down_tlast),
    .up_xfcp_in_tuser(xfcp_qsfp2_gty_down_tuser),
    .up_xfcp_out_tdata(xfcp_qsfp2_gty_up_tdata),
    .up_xfcp_out_tvalid(xfcp_qsfp2_gty_up_tvalid),
    .up_xfcp_out_tready(xfcp_qsfp2_gty_up_tready),
    .up_xfcp_out_tlast(xfcp_qsfp2_gty_up_tlast),
    .up_xfcp_out_tuser(xfcp_qsfp2_gty_up_tuser),

    .gty_com_drp_addr(qsfp_gty_com_drp_addr[1*10 +: 10]),
    .gty_com_drp_do(qsfp_gty_com_drp_do[1*16 +: 16]),
    .gty_com_drp_di(qsfp_gty_com_drp_di[1*16 +: 16]),
    .gty_com_drp_en(qsfp_gty_com_drp_en[1*1 +: 1]),
    .gty_com_drp_we(qsfp_gty_com_drp_we[1*1 +: 1]),
    .gty_com_drp_rdy(qsfp_gty_com_drp_rdy[1*1 +: 1]),

    .gty_drp_addr(qsfp_gty_drp_addr[1*4*10 +: 4*10]),
    .gty_drp_do(qsfp_gty_drp_do[1*4*16 +: 4*16]),
    .gty_drp_di(qsfp_gty_drp_di[1*4*16 +: 4*16]),
    .gty_drp_en(qsfp_gty_drp_en[1*4*1 +: 4*1]),
    .gty_drp_we(qsfp_gty_drp_we[1*4*1 +: 4*1]),
    .gty_drp_rdy(qsfp_gty_drp_rdy[1*4*1 +: 4*1]),

    .gty_reset(qsfp_gty_reset[1*4*1 +: 4*1]),
    .gty_tx_reset(qsfp_gty_tx_reset[1*4*1 +: 4*1]),
    .gty_rx_reset(qsfp_gty_rx_reset[1*4*1 +: 4*1]),

    .gty_txusrclk2({4{qsfp_gty_txusrclk2}}),
    .gty_txprbssel(qsfp_gty_txprbssel[1*4*4 +: 4*4]),
    .gty_txprbsforceerr(qsfp_gty_txprbsforceerr[1*4*1 +: 4*1]),
    .gty_txpolarity(qsfp_gty_txpolarity[1*4*1 +: 4*1]),
    .gty_txelecidle(qsfp_gty_txelecidle[1*4*1 +: 4*1]),
    .gty_txinhibit(qsfp_gty_txinhibit[1*4*1 +: 4*1]),
    .gty_txdiffctrl(qsfp_gty_txdiffctrl[1*4*5 +: 4*5]),
    .gty_txmaincursor(qsfp_gty_txmaincursor[1*4*7 +: 4*7]),
    .gty_txpostcursor(qsfp_gty_txpostcursor[1*4*5 +: 4*5]),
    .gty_txprecursor(qsfp_gty_txprecursor[1*4*5 +: 4*5]),

    .gty_rxusrclk2({4{qsfp_gty_rxusrclk2}}),
    .gty_rxpolarity(qsfp_gty_rxpolarity[1*4*1 +: 4*1]),
    .gty_rxprbscntreset(qsfp_gty_rxprbscntreset[1*4*1 +: 4*1]),
    .gty_rxprbssel(qsfp_gty_rxprbssel[1*4*4 +: 4*4]),
    .gty_rxprbserr(qsfp_gty_rxprbserr[1*4*1 +: 4*1]),
    .gty_rxprbslocked(qsfp_gty_rxprbslocked[1*4*1 +: 4*1])
);

wire qsfp1_mgt_refclk_0;

IBUFDS_GTE4 ibufds_gte4_qsfp1_mgt_refclk_0_inst (
    .I             (qsfp1_mgt_refclk_0_p),
    .IB            (qsfp1_mgt_refclk_0_n),
    .CEB           (1'b0),
    .O             (qsfp1_mgt_refclk_0),
    .ODIV2         ()
);

gtwizard_ultrascale_0 gtwizard_ultrascale_0_inst (
    .gtyrxn_in                           ({qsfp2_rx4_n, qsfp2_rx3_n, qsfp2_rx2_n, qsfp2_rx1_n, qsfp1_rx4_n, qsfp1_rx3_n, qsfp1_rx2_n, qsfp1_rx1_n}),
    .gtyrxp_in                           ({qsfp2_rx4_p, qsfp2_rx3_p, qsfp2_rx2_p, qsfp2_rx1_p, qsfp1_rx4_p, qsfp1_rx3_p, qsfp1_rx2_p, qsfp1_rx1_p}),
    .gtytxn_out                          ({qsfp2_tx4_n, qsfp2_tx3_n, qsfp2_tx2_n, qsfp2_tx1_n, qsfp1_tx4_n, qsfp1_tx3_n, qsfp1_tx2_n, qsfp1_tx1_n}),
    .gtytxp_out                          ({qsfp2_tx4_p, qsfp2_tx3_p, qsfp2_tx2_p, qsfp2_tx1_p, qsfp1_tx4_p, qsfp1_tx3_p, qsfp1_tx2_p, qsfp1_tx1_p}),
    .gtwiz_userclk_tx_reset_in           (gty_drp_rst),
    .gtwiz_userclk_tx_srcclk_out         (),
    .gtwiz_userclk_tx_usrclk_out         (),
    .gtwiz_userclk_tx_usrclk2_out        (qsfp_gty_txusrclk2),
    .gtwiz_userclk_tx_active_out         (),
    .gtwiz_userclk_rx_reset_in           (gty_drp_rst),
    .gtwiz_userclk_rx_srcclk_out         (),
    .gtwiz_userclk_rx_usrclk_out         (),
    .gtwiz_userclk_rx_usrclk2_out        (qsfp_gty_rxusrclk2),
    .gtwiz_userclk_rx_active_out         (),
    .gtwiz_reset_clk_freerun_in          (gty_drp_clk),
    .gtwiz_reset_all_in                  (gty_drp_rst || qsfp_gty_reset),
    .gtwiz_reset_tx_pll_and_datapath_in  (|qsfp_gty_tx_reset),
    .gtwiz_reset_tx_datapath_in          (1'b0),
    .gtwiz_reset_rx_pll_and_datapath_in  (|qsfp_gty_rx_reset),
    .gtwiz_reset_rx_datapath_in          (1'b0),
    .gtwiz_reset_rx_cdr_stable_out       (),
    .gtwiz_reset_tx_done_out             (),
    .gtwiz_reset_rx_done_out             (),
    .gtwiz_userdata_tx_in                ({8{64'd0}}),
    .gtwiz_userdata_rx_out               (),
    .drpaddr_common_in                   (qsfp_gty_com_drp_addr),
    .drpclk_common_in                    ({2{gty_drp_clk}}),
    .drpdi_common_in                     (qsfp_gty_com_drp_do),
    .drpen_common_in                     (qsfp_gty_com_drp_en),
    .drpwe_common_in                     (qsfp_gty_com_drp_we),
    .gtrefclk00_in                       ({2{qsfp1_mgt_refclk_0}}),
    .drpdo_common_out                    (qsfp_gty_com_drp_di),
    .drprdy_common_out                   (qsfp_gty_com_drp_rdy),
    .qpll0outclk_out                     (),
    .qpll0outrefclk_out                  (),
    .drpaddr_in                          (qsfp_gty_drp_addr),
    .drpclk_in                           ({8{gty_drp_clk}}),
    .drpdi_in                            (qsfp_gty_drp_do),
    .drpen_in                            (qsfp_gty_drp_en),
    .drpwe_in                            (qsfp_gty_drp_we),
    .rxpolarity_in                       (qsfp_gty_rxpolarity),
    .rxprbscntreset_in                   (qsfp_gty_rxprbscntreset),
    .rxprbssel_in                        (qsfp_gty_rxprbssel),
    .txdiffctrl_in                       (qsfp_gty_txdiffctrl),
    .txelecidle_in                       (qsfp_gty_txelecidle),
    .txinhibit_in                        (qsfp_gty_txinhibit),
    .txmaincursor_in                     (qsfp_gty_txmaincursor),
    .txpolarity_in                       (qsfp_gty_txpolarity),
    .txpostcursor_in                     (qsfp_gty_txpostcursor),
    .txprbsforceerr_in                   (qsfp_gty_txprbsforceerr),
    .txprbssel_in                        (qsfp_gty_txprbssel),
    .txprecursor_in                      (qsfp_gty_txprecursor),
    .drpdo_out                           (qsfp_gty_drp_di),
    .drprdy_out                          (qsfp_gty_drp_rdy),
    .rxpmaresetdone_out                  (),
    .rxprbserr_out                       (qsfp_gty_rxprbserr),
    .rxprbslocked_out                    (qsfp_gty_rxprbslocked),
    .txpmaresetdone_out                  (),
    .txprgdivresetdone_out               ()
);

// SGMII interface to PHY
wire phy_gmii_clk_int;
wire phy_gmii_rst_int;
wire phy_gmii_clk_en_int;
wire [7:0] phy_gmii_txd_int;
wire phy_gmii_tx_en_int;
wire phy_gmii_tx_er_int;
wire [7:0] phy_gmii_rxd_int;
wire phy_gmii_rx_dv_int;
wire phy_gmii_rx_er_int;

wire [15:0] gig_eth_pcspma_status_vector;

wire gig_eth_pcspma_status_link_status              = gig_eth_pcspma_status_vector[0];
wire gig_eth_pcspma_status_link_synchronization     = gig_eth_pcspma_status_vector[1];
wire gig_eth_pcspma_status_rudi_c                   = gig_eth_pcspma_status_vector[2];
wire gig_eth_pcspma_status_rudi_i                   = gig_eth_pcspma_status_vector[3];
wire gig_eth_pcspma_status_rudi_invalid             = gig_eth_pcspma_status_vector[4];
wire gig_eth_pcspma_status_rxdisperr                = gig_eth_pcspma_status_vector[5];
wire gig_eth_pcspma_status_rxnotintable             = gig_eth_pcspma_status_vector[6];
wire gig_eth_pcspma_status_phy_link_status          = gig_eth_pcspma_status_vector[7];
wire [1:0] gig_eth_pcspma_status_remote_fault_encdg = gig_eth_pcspma_status_vector[9:8];
wire [1:0] gig_eth_pcspma_status_speed              = gig_eth_pcspma_status_vector[11:10];
wire gig_eth_pcspma_status_duplex                   = gig_eth_pcspma_status_vector[12];
wire gig_eth_pcspma_status_remote_fault             = gig_eth_pcspma_status_vector[13];
wire [1:0] gig_eth_pcspma_status_pause              = gig_eth_pcspma_status_vector[15:14];

wire [4:0] gig_eth_pcspma_config_vector;

assign gig_eth_pcspma_config_vector[4] = 1'b1; // autonegotiation enable
assign gig_eth_pcspma_config_vector[3] = 1'b0; // isolate
assign gig_eth_pcspma_config_vector[2] = 1'b0; // power down
assign gig_eth_pcspma_config_vector[1] = 1'b0; // loopback enable
assign gig_eth_pcspma_config_vector[0] = 1'b0; // unidirectional enable

wire [15:0] gig_eth_pcspma_an_config_vector;

assign gig_eth_pcspma_an_config_vector[15]    = 1'b1;    // SGMII link status
assign gig_eth_pcspma_an_config_vector[14]    = 1'b1;    // SGMII Acknowledge
assign gig_eth_pcspma_an_config_vector[13:12] = 2'b01;   // full duplex
assign gig_eth_pcspma_an_config_vector[11:10] = 2'b10;   // SGMII speed
assign gig_eth_pcspma_an_config_vector[9]     = 1'b0;    // reserved
assign gig_eth_pcspma_an_config_vector[8:7]   = 2'b00;   // pause frames - SGMII reserved
assign gig_eth_pcspma_an_config_vector[6]     = 1'b0;    // reserved
assign gig_eth_pcspma_an_config_vector[5]     = 1'b0;    // full duplex - SGMII reserved
assign gig_eth_pcspma_an_config_vector[4:1]   = 4'b0000; // reserved
assign gig_eth_pcspma_an_config_vector[0]     = 1'b1;    // SGMII

gig_ethernet_pcs_pma_0 
eth_pcspma (
    // SGMII
    .txp_0                  (phy_sgmii_tx_p),
    .txn_0                  (phy_sgmii_tx_n),
    .rxp_0                  (phy_sgmii_rx_p),
    .rxn_0                  (phy_sgmii_rx_n),

    // Ref clock from PHY
    .refclk625_p            (phy_sgmii_clk_p),
    .refclk625_n            (phy_sgmii_clk_n),

    // async reset
    .reset                  (rst_125mhz_int),

    // clock and reset outputs
    .clk125_out             (phy_gmii_clk_int),
    .clk312_out             (),
    .rst_125_out            (phy_gmii_rst_int),
    .tx_logic_reset         (),
    .rx_logic_reset         (),
    .tx_locked              (),
    .rx_locked              (),
    .tx_pll_clk_out         (),
    .rx_pll_clk_out         (),

    // MAC clocking
    .sgmii_clk_r_0          (),
    .sgmii_clk_f_0          (),
    .sgmii_clk_en_0         (phy_gmii_clk_en_int),
    
    // Speed control
    .speed_is_10_100_0      (gig_eth_pcspma_status_speed != 2'b10),
    .speed_is_100_0         (gig_eth_pcspma_status_speed == 2'b01),

    // Internal GMII
    .gmii_txd_0             (phy_gmii_txd_int),
    .gmii_tx_en_0           (phy_gmii_tx_en_int),
    .gmii_tx_er_0           (phy_gmii_tx_er_int),
    .gmii_rxd_0             (phy_gmii_rxd_int),
    .gmii_rx_dv_0           (phy_gmii_rx_dv_int),
    .gmii_rx_er_0           (phy_gmii_rx_er_int),
    .gmii_isolate_0         (),

    // Configuration
    .configuration_vector_0 (gig_eth_pcspma_config_vector),

    .an_interrupt_0         (),
    .an_adv_config_vector_0 (gig_eth_pcspma_an_config_vector),
    .an_restart_config_0    (1'b0),

    // Status
    .status_vector_0        (gig_eth_pcspma_status_vector),
    .signal_detect_0        (1'b1),

    // Cascade
    .tx_bsc_rst_out         (),
    .rx_bsc_rst_out         (),
    .tx_bs_rst_out          (),
    .rx_bs_rst_out          (),
    .tx_rst_dly_out         (),
    .rx_rst_dly_out         (),
    .tx_bsc_en_vtc_out      (),
    .rx_bsc_en_vtc_out      (),
    .tx_bs_en_vtc_out       (),
    .rx_bs_en_vtc_out       (),
    .riu_clk_out            (),
    .riu_addr_out           (),
    .riu_wr_data_out        (),
    .riu_wr_en_out          (),
    .riu_nibble_sel_out     (),
    .riu_rddata_1           (16'b0),
    .riu_valid_1            (1'b0),
    .riu_prsnt_1            (1'b0),
    .riu_rddata_2           (16'b0),
    .riu_valid_2            (1'b0),
    .riu_prsnt_2            (1'b0),
    .riu_rddata_3           (16'b0),
    .riu_valid_3            (1'b0),
    .riu_prsnt_3            (1'b0),
    .rx_btval_1             (),
    .rx_btval_2             (),
    .rx_btval_3             (),
    .tx_dly_rdy_1           (1'b1),
    .rx_dly_rdy_1           (1'b1),
    .rx_vtc_rdy_1           (1'b1),
    .tx_vtc_rdy_1           (1'b1),
    .tx_dly_rdy_2           (1'b1),
    .rx_dly_rdy_2           (1'b1),
    .rx_vtc_rdy_2           (1'b1),
    .tx_vtc_rdy_2           (1'b1),
    .tx_dly_rdy_3           (1'b1),
    .rx_dly_rdy_3           (1'b1),
    .rx_vtc_rdy_3           (1'b1),
    .tx_vtc_rdy_3           (1'b1),
    .tx_rdclk_out           ()
);

reg [19:0] delay_reg = 20'hfffff;

reg [4:0] mdio_cmd_phy_addr = 5'h03;
reg [4:0] mdio_cmd_reg_addr = 5'h00;
reg [15:0] mdio_cmd_data = 16'd0;
reg [1:0] mdio_cmd_opcode = 2'b01;
reg mdio_cmd_valid = 1'b0;
wire mdio_cmd_ready;

reg [3:0] state_reg = 0;

always @(posedge clk_125mhz_int) begin
    if (rst_125mhz_int) begin
        state_reg <= 0;
        delay_reg <= 20'hfffff;
        mdio_cmd_reg_addr <= 5'h00;
        mdio_cmd_data <= 16'd0;
        mdio_cmd_valid <= 1'b0;
    end else begin
        mdio_cmd_valid <= mdio_cmd_valid & !mdio_cmd_ready;
        if (delay_reg > 0) begin
            delay_reg <= delay_reg - 1;
        end else if (!mdio_cmd_ready) begin
            // wait for ready
            state_reg <= state_reg;
        end else begin
            mdio_cmd_valid <= 1'b0;
            case (state_reg)
                // set SGMII autonegotiation timer to 11 ms
                // write 0x0070 to CFG4 (0x0031)
                4'd0: begin
                    // write to REGCR to load address
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h001F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd1;
                end
                4'd1: begin
                    // write address of CFG4 to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h0031;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd2;
                end
                4'd2: begin
                    // write to REGCR to load data
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h401F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd3;
                end
                4'd3: begin
                    // write data for CFG4 to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h0070;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd4;
                end
                // enable SGMII clock output
                // write 0x4000 to SGMIICTL1 (0x00D3)
                4'd4: begin
                    // write to REGCR to load address
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h001F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd5;
                end
                4'd5: begin
                    // write address of SGMIICTL1 to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h00D3;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd6;
                end
                4'd6: begin
                    // write to REGCR to load data
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h401F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd7;
                end
                4'd7: begin
                    // write data for SGMIICTL1 to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h4000;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd8;
                end
                // enable 10Mbps operation
                // write 0x0015 to 10M_SGMII_CFG (0x016F)
                4'd8: begin
                    // write to REGCR to load address
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h001F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd9;
                end
                4'd9: begin
                    // write address of 10M_SGMII_CFG to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h016F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd10;
                end
                4'd10: begin
                    // write to REGCR to load data
                    mdio_cmd_reg_addr <= 5'h0D;
                    mdio_cmd_data <= 16'h401F;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd11;
                end
                4'd11: begin
                    // write data for 10M_SGMII_CFG to ADDAR
                    mdio_cmd_reg_addr <= 5'h0E;
                    mdio_cmd_data <= 16'h0015;
                    mdio_cmd_valid <= 1'b1;
                    state_reg <= 4'd12;
                end
                4'd12: begin
                    // done
                    state_reg <= 4'd12;
                end
            endcase
        end
    end
end

wire mdc;
wire mdio_i;
wire mdio_o;
wire mdio_t;

mdio_master
mdio_master_inst (
    .clk(clk_125mhz_int),
    .rst(rst_125mhz_int),

    .cmd_phy_addr(mdio_cmd_phy_addr),
    .cmd_reg_addr(mdio_cmd_reg_addr),
    .cmd_data(mdio_cmd_data),
    .cmd_opcode(mdio_cmd_opcode),
    .cmd_valid(mdio_cmd_valid),
    .cmd_ready(mdio_cmd_ready),

    .data_out(),
    .data_out_valid(),
    .data_out_ready(1'b1),

    .mdc_o(mdc),
    .mdio_i(mdio_i),
    .mdio_o(mdio_o),
    .mdio_t(mdio_t),

    .busy(),

    .prescale(8'd3)
);

assign phy_mdc = mdc;
assign mdio_i = phy_mdio;
assign phy_mdio = mdio_t ? 1'bz : mdio_o;

fpga_core
core_inst (
    /*
     * Clock: 125MHz
     * Synchronous reset
     */
    .clk(clk_125mhz_int),
    .rst(rst_125mhz_int),
    /*
     * GPIO
     */
    .btnu(btnu_int),
    .btnl(btnl_int),
    .btnd(btnd_int),
    .btnr(btnr_int),
    .btnc(btnc_int),
    .sw(sw_int),
    .led(led),
    /*
     * I2C
     */
    .i2c_scl_i(i2c_scl_i),
    .i2c_scl_o(i2c_scl_o),
    .i2c_scl_t(i2c_scl_t),
    .i2c_sda_i(i2c_sda_i),
    .i2c_sda_o(i2c_sda_o),
    .i2c_sda_t(i2c_sda_t),
    /*
     * Ethernet: 1000BASE-T SGMII
     */
    .phy_gmii_clk(phy_gmii_clk_int),
    .phy_gmii_rst(phy_gmii_rst_int),
    .phy_gmii_clk_en(phy_gmii_clk_en_int),
    .phy_gmii_rxd(phy_gmii_rxd_int),
    .phy_gmii_rx_dv(phy_gmii_rx_dv_int),
    .phy_gmii_rx_er(phy_gmii_rx_er_int),
    .phy_gmii_txd(phy_gmii_txd_int),
    .phy_gmii_tx_en(phy_gmii_tx_en_int),
    .phy_gmii_tx_er(phy_gmii_tx_er_int),
    .phy_reset_n(phy_reset_n),
    .phy_int_n(phy_int_n),
    /*
     * UART: 115200 bps, 8N1
     */
    .uart_rxd(uart_rxd_int),
    .uart_txd(uart_txd),
    .uart_rts(uart_rts),
    .uart_cts(uart_cts_int),
    /*
     * Transceiver control
     */
    .xfcp_mgt_up_tdata(xfcp_mgt_up_tdata),
    .xfcp_mgt_up_tvalid(xfcp_mgt_up_tvalid),
    .xfcp_mgt_up_tready(xfcp_mgt_up_tready),
    .xfcp_mgt_up_tlast(xfcp_mgt_up_tlast),
    .xfcp_mgt_up_tuser(xfcp_mgt_up_tuser),
    .xfcp_mgt_down_tdata(xfcp_mgt_down_tdata),
    .xfcp_mgt_down_tvalid(xfcp_mgt_down_tvalid),
    .xfcp_mgt_down_tready(xfcp_mgt_down_tready),
    .xfcp_mgt_down_tlast(xfcp_mgt_down_tlast),
    .xfcp_mgt_down_tuser(xfcp_mgt_down_tuser)
);

endmodule
